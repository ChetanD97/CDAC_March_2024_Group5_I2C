module tb;
   
